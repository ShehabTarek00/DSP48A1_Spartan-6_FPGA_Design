module Main_DSP_TB();
reg [17:0]A_TB,B_TB,BCIN_TB,D_TB;
reg [47:0]C_TB,PCIN_TB;

reg[7:0]opmode_TB;
reg CARRYIN_TB;
wire [47:0]P_DUT;
wire CARRYOUT_DUT;
reg [47:0]P_EXP;
reg CARRYOUT_EXP;
wire [35:0]M_DUT;
reg [35:0]M_EXP;
wire [17:0]BCOUT_DUT;
reg [17:0]BCOUT_EXP;
wire CARRYOUTF_DUT;
reg CARRYOUTF_EXP;

wire [47:0]PCOUT_DUT;
reg [47:0]PCOUT_EXP;

reg [47:0]buffer;
reg CLK_TB,CEA_TB,CEB_TB,CEC_TB,CECARRYIN_TB,CED_TB,CEM_TB,
CEOPMODE_TB,CEP_TB,
RSTA_TB,RSTB_TB,RSTC_TB,RSTCARRYIN_TB,
RSTD_TB,RSTM_TB,RSTOPMODE_TB,RSTP_TB;


Main_DSP DUT(A_TB,B_TB,C_TB,D_TB,CARRYIN_TB,M_DUT,P_DUT,
	CARRYOUT_DUT,CARRYOUTF_DUT,CLK_TB,opmode_TB,
CEA_TB,CEB_TB,CEC_TB,CECARRYIN_TB,CED_TB,CEM_TB,CEOPMODE_TB,CEP_TB,
RSTA_TB,RSTB_TB,RSTC_TB,RSTCARRYIN_TB,RSTD_TB,RSTM_TB,RSTOPMODE_TB,
RSTP_TB,BCIN_TB,BCOUT_DUT,PCOUT_DUT,PCIN_TB);


initial begin
	CLK_TB=0;
	forever 
	#1 CLK_TB=~CLK_TB;
end

initial begin
	#0 
CEA_TB=1;CEB_TB=1;CEC_TB=1;CED_TB=1;
	CECARRYIN_TB=1;CEOPMODE_TB=1;CEM_TB=1;CEP_TB=1;

RSTA_TB=0;RSTB_TB=0;RSTC_TB=0;RSTCARRYIN_TB=0;RSTD_TB=0;
RSTM_TB=0;RSTOPMODE_TB=0;RSTP_TB=0;

A_TB=18'hA7; B_TB=18'hB7; C_TB=48'hC7; D_TB=18'hD7;
opmode_TB=8'b0_0_0_1_11_01;PCIN_TB=$random;BCIN_TB=$random;
CARRYIN_TB=$random;
BCOUT_EXP=18'h18E;M_EXP=36'h103A2;
#7
PCOUT_EXP=48'h10469;P_EXP=48'h10469;
CARRYOUT_EXP=0;CARRYOUTF_EXP=0;
#20
if ((BCOUT_EXP != BCOUT_DUT) || (M_EXP != M_DUT) || (PCOUT_DUT != PCOUT_EXP) || (P_DUT != P_EXP) || (CARRYOUT_DUT != CARRYOUT_EXP) || (CARRYOUTF_DUT != CARRYOUTF_EXP)) begin
	$display("Error here");
	$stop;
end



	#20 
CEA_TB=1;CEB_TB=1;CEC_TB=1;CED_TB=1;
	CECARRYIN_TB=1;CEOPMODE_TB=1;CEM_TB=1;CEP_TB=1;

RSTA_TB=1;RSTB_TB=1;RSTC_TB=1;RSTCARRYIN_TB=1;RSTD_TB=1;
RSTM_TB=1;RSTOPMODE_TB=1;RSTP_TB=1;

A_TB=18'hA7; B_TB=18'hB7; C_TB=48'hC7; D_TB=18'hD7;
opmode_TB=8'b0_0_0_1_11_01;PCIN_TB=$random;BCIN_TB=$random;
CARRYIN_TB=$random;
BCOUT_EXP=18'h0;M_EXP=36'h0;
#7
PCOUT_EXP=48'h0;P_EXP=48'h0;
CARRYOUT_EXP=0;CARRYOUTF_EXP=0;
#20
if ((BCOUT_EXP != BCOUT_DUT) || (M_EXP != M_DUT) || (PCOUT_DUT != PCOUT_EXP) || (P_DUT != P_EXP) || (CARRYOUT_DUT != CARRYOUT_EXP) || (CARRYOUTF_DUT != CARRYOUTF_EXP)) begin
	$display("Error here");
	$stop;
end

#20 
CEA_TB=1;CEB_TB=1;CEC_TB=1;CED_TB=1;
	CECARRYIN_TB=1;CEOPMODE_TB=1;CEM_TB=1;CEP_TB=1;

RSTA_TB=0;RSTB_TB=0;RSTC_TB=0;RSTCARRYIN_TB=0;RSTD_TB=0;
RSTM_TB=0;RSTOPMODE_TB=0;RSTP_TB=0;

A_TB=18'hA7; B_TB=18'hB7; C_TB=48'hCCC7; D_TB=18'hD7;
opmode_TB=8'b1_1_1_1_11_01;PCIN_TB=$random;BCIN_TB=$random;
CARRYIN_TB=$random;
BCOUT_EXP=18'h20;M_EXP=36'h14E0;
#7
PCOUT_EXP=48'hB7E6;P_EXP=48'hB7E6;
CARRYOUT_EXP=0;CARRYOUTF_EXP=0;
#20
if ((BCOUT_EXP != BCOUT_DUT) || (M_EXP != M_DUT) || (PCOUT_DUT != PCOUT_EXP) || (P_DUT != P_EXP) || (CARRYOUT_DUT != CARRYOUT_EXP) || (CARRYOUTF_DUT != CARRYOUTF_EXP)) begin
	$display("Error here");
	$stop;
end


#20 
CEA_TB=1;CEB_TB=1;CEC_TB=1;CED_TB=1;
	CECARRYIN_TB=1;CEOPMODE_TB=1;CEM_TB=1;CEP_TB=1;

RSTA_TB=0;RSTB_TB=0;RSTC_TB=0;RSTCARRYIN_TB=0;RSTD_TB=0;
RSTM_TB=0;RSTOPMODE_TB=0;RSTP_TB=0;

A_TB=18'hA7; B_TB=18'hB7; C_TB=48'hCCC7; D_TB=18'hD7;
opmode_TB=8'b0_0_0_0_01_01;PCIN_TB=48'h1221;BCIN_TB=$random;
CARRYIN_TB=$random;
BCOUT_EXP=18'hB7;M_EXP=36'h7761;
#7
PCOUT_EXP=48'h8982;P_EXP=48'h8982;
CARRYOUT_EXP=0;CARRYOUTF_EXP=0;
#20
if ((BCOUT_EXP != BCOUT_DUT) || (M_EXP != M_DUT) || (PCOUT_DUT != PCOUT_EXP) || (P_DUT != P_EXP) || (CARRYOUT_DUT != CARRYOUT_EXP) || (CARRYOUTF_DUT != CARRYOUTF_EXP)) begin
	$display("Error here");
	$stop;
end
buffer=PCOUT_EXP;
#20 
CEA_TB=1;CEB_TB=1;CEC_TB=1;CED_TB=1;
	CECARRYIN_TB=1;CEOPMODE_TB=1;CEM_TB=1;CEP_TB=1;

RSTA_TB=0;RSTB_TB=0;RSTC_TB=0;RSTCARRYIN_TB=0;RSTD_TB=0;
RSTM_TB=0;RSTOPMODE_TB=0;RSTP_TB=0;

A_TB=18'hA7; B_TB=18'hB7; C_TB=48'hCCC7; D_TB=18'hD7;
opmode_TB=8'b0_0_0_1_10_00;PCIN_TB=48'h1221;BCIN_TB=$random;
CARRYIN_TB=$random;
BCOUT_EXP=18'h18E;M_EXP=36'h103A2;
#7
PCOUT_EXP=buffer;P_EXP=buffer;
CARRYOUT_EXP=0;CARRYOUTF_EXP=0;
#20
if ((BCOUT_EXP != BCOUT_DUT) || (M_EXP != M_DUT) || (PCOUT_DUT != PCOUT_EXP) || (P_DUT != P_EXP) || (CARRYOUT_DUT != CARRYOUT_EXP) || (CARRYOUTF_DUT != CARRYOUTF_EXP)) begin
	$display("Error here");
	$stop;
end


#20 
CEA_TB=1;CEB_TB=1;CEC_TB=1;CED_TB=1;
	CECARRYIN_TB=1;CEOPMODE_TB=1;CEM_TB=1;CEP_TB=1;

RSTA_TB=0;RSTB_TB=0;RSTC_TB=0;RSTCARRYIN_TB=0;RSTD_TB=0;
RSTM_TB=0;RSTOPMODE_TB=0;RSTP_TB=0;

A_TB=18'h3FFFF; B_TB=18'hB; C_TB=48'hCCC7; D_TB=18'hD;
opmode_TB=8'b0_0_0_1_00_11;PCIN_TB=48'h1221;BCIN_TB=$random;
CARRYIN_TB=$random;
BCOUT_EXP=18'h18;M_EXP=36'h5FFFE8;
#7
PCOUT_EXP=48'hDFFFFC0018;P_EXP=48'hDFFFFC0018;
CARRYOUT_EXP=0;CARRYOUTF_EXP=0;
#20
if ((BCOUT_EXP != BCOUT_DUT) || (M_EXP != M_DUT) || (PCOUT_DUT != PCOUT_EXP) || (P_DUT != P_EXP) || (CARRYOUT_DUT != CARRYOUT_EXP) || (CARRYOUTF_DUT != CARRYOUTF_EXP)) begin
	$display("Error here");
	$stop;
end



end//of the main initial

initial begin
	$monitor("A=%h,B=%h,C=%h,D=%h,M=%h,BCOUT=%h,P=%h",A_TB,B_TB,C_TB,D_TB,M_EXP,BCOUT_EXP,P_EXP);
end
endmodule